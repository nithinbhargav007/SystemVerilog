
//calendar scheduling for 3 people ( 5 days of the week, 90 mins slot each)

module calendar_scheduling;
  initial begin
    
    string person1[string][string] = { "Monday":'{"0000":"No","0130":"No","0300":"Yes","0430":"No","0600":"Yes","0730":"Yes","0900":"No",
                                       "1030":"Yes","1200":"No","1330":"Yes","1500":"No","1630":"Yes","1800":"Yes","1930":"No","21:00":"Yes","2230":"Yes"},
                                        "Tuesday":'{"0000":"Yes","0130":"No","0300":"Yes","0430":"No","0600":"Yes","0730":"Yes","0900":"No",
                                       "1030":"Yes","1200":"No","1330":"Yes","1500":"No","1630":"Yes","1800":"Yes","1930":"No","21:00":"Yes","2230":"Yes"},
                                        "Wednesday":'{"0000":"Yes","0130":"No","0300":"Yes","0430":"No","0600":"Yes","0730":"Yes","0900":"No",
                                       "1030":"Yes","1200":"No","1330":"Yes","1500":"No","1630":"Yes","1800":"Yes","1930":"No","21:00":"Yes","2230":"Yes"},
                                        "Thursday":'{"0000":"Yes","0130":"No","0300":"Yes","0430":"No","0600":"Yes","0730":"Yes","0900":"No",
                                       "1030":"Yes","1200":"No","1330":"Yes","1500":"No","1630":"Yes","1800":"Yes","1930":"No","21:00":"Yes","2230":"Yes"},
                                        "Friday":'{"0000":"Yes","0130":"No","0300":"Yes","0430":"No","0600":"Yes","0730":"Yes","0900":"No",
                                       "1030":"Yes","1200":"No","1330":"Yes","1500":"No","1630":"Yes","1800":"Yes","1930":"No","21:00":"Yes","2230":"Yes"}
                                       };
                             
    string person2[string][string] = {"Monday":'{"0000":"No","0130":"Yes","0300":"No","0430":"Yes","0600":"Yes","0730":"Yes","0900":"No",
                                      "1030":"No","1200":"No","1330":"No","1500":"No","1630":"Yes","1800":"No","1930":"Yes","21:00":"No","2230":"Yes"},
                                      "Tuesday":'{"0000":"Yes","0130":"Yes","0300":"No","0430":"Yes","0600":"Yes","0730":"Yes","0900":"No",
                                      "1030":"No","1200":"No","1330":"No","1500":"No","1630":"Yes","1800":"No","1930":"Yes","21:00":"No","2230":"Yes"},
                                      "Wednesday":'{"0000":"Yes","0130":"Yes","0300":"No","0430":"Yes","0600":"Yes","0730":"Yes","0900":"No",
                                      "1030":"No","1200":"No","1330":"No","1500":"No","1630":"Yes","1800":"No","1930":"Yes","21:00":"No","2230":"Yes"},
                                      "Thursday":'{"0000":"Yes","0130":"Yes","0300":"No","0430":"Yes","0600":"Yes","0730":"Yes","0900":"No",
                                      "1030":"No","1200":"No","1330":"No","1500":"No","1630":"Yes","1800":"No","1930":"Yes","21:00":"No","2230":"Yes"},
                                      "Friday":'{"0000":"Yes","0130":"Yes","0300":"No","0430":"Yes","0600":"Yes","0730":"Yes","0900":"No",
                                      "1030":"No","1200":"No","1330":"No","1500":"No","1630":"Yes","1800":"No","1930":"Yes","21:00":"No","2230":"Yes"}
                                     };
  
    string person3[string][string] = {"Monday":'{"0000":"No","0130":"Yes","0300":"Yes","0430":"Yes","0600":"Yes","0730":"Yes","0900":"Yes",
                                       "1030":"Yes","1200":"No","1330":"Yes","1500":"No","1630":"No","1800":"No","1930":"No","21:00":"No","2230":"Yes"},
                                      "Tuesday":'{"0000":"Yes","0130":"Yes","0300":"Yes","0430":"Yes","0600":"Yes","0730":"Yes","0900":"Yes",
                                       "1030":"Yes","1200":"No","1330":"Yes","1500":"No","1630":"No","1800":"No","1930":"No","21:00":"No","2230":"Yes"},
                                      "Wednesday":'{"0000":"Yes","0130":"Yes","0300":"Yes","0430":"Yes","0600":"Yes","0730":"Yes","0900":"Yes",
                                       "1030":"Yes","1200":"No","1330":"Yes","1500":"No","1630":"No","1800":"No","1930":"No","21:00":"No","2230":"Yes"},
                                       "Thursday":'{"0000":"Yes","0130":"Yes","0300":"Yes","0430":"Yes","0600":"Yes","0730":"Yes","0900":"Yes",
                                       "1030":"Yes","1200":"No","1330":"Yes","1500":"No","1630":"No","1800":"No","1930":"No","21:00":"No","2230":"Yes"},
                                        "Friday":'{"0000":"Yes","0130":"Yes","0300":"Yes","0430":"Yes","0600":"Yes","0730":"Yes","0900":"Yes",
                                       "1030":"Yes","1200":"No","1330":"Yes","1500":"No","1630":"No","1800":"No","1930":"No","21:00":"No","2230":"Yes"}
    								 };

    foreach(person1[i,j]) begin
      //$display("The calendar values are as follows Time : %0s :  %0s  : %0s : %0s : %0s",i,j,person1[i][j],person2[i][j],person3[i][j]);
      if((person1[i][j]==person2[i][j])&&(person2[i][j]==person3[i][j]))
        $display("All the three people are available at time %0s IST on %0s", j, i);
    end    
  end
  
endmodule